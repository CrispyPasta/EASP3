module ALU( data_in, operation, data_out);

input data_in;
input operation;
output data_out;

assign data_out = data_in;


endmodule