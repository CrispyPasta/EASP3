module Memory(MAR_value, data_input, MBR_value, clk);

input [7:0] MAR_value;
input [7:0] data_input;
output [7:0] MBR_value;
input clk;


endmodule