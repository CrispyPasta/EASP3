module Prac3();

Memory my_Memory(MAR_value, data_input, MBR_value, clk);
CPU my_CPU( MAR_value, MBR_value, clk );

endmodule